library verilog;
use verilog.vl_types.all;
entity lab2_if is
    port(
        clk             : in     vl_logic
    );
end lab2_if;
